module dbg_bridge_fifo
//-----------------------------------------------------------------
// Params
//-----------------------------------------------------------------
#(
    parameter WIDTH  = 8,
    parameter DEPTH  = 4,
    parameter ADDR_W = 2
)
//-----------------------------------------------------------------
// Ports
//-----------------------------------------------------------------
(
    // Inputs
    input             clk_i,
    input             rst_i,
    input [WIDTH-1:0] data_in_i,
    input             push_i,
    input             pop_i,

    // Outputs
    output [WIDTH-1:0] data_out_o,
    output             accept_o,
    output             valid_o
);

  //-----------------------------------------------------------------
  // Local Params
  //-----------------------------------------------------------------
  localparam COUNT_W = ADDR_W + 1;

  //-----------------------------------------------------------------
  // Registers
  //-----------------------------------------------------------------
  reg [WIDTH-1:0] ram_q[DEPTH-1:0];
  reg [ADDR_W-1:0] rd_ptr_q;
  reg [ADDR_W-1:0] wr_ptr_q;
  reg [COUNT_W-1:0] count_q;

  //-----------------------------------------------------------------
  // Sequential
  //-----------------------------------------------------------------
  always @(posedge clk_i or negedge rst_i)
    if (!rst_i) begin
      count_q  <= {(COUNT_W) {1'b0}};
      rd_ptr_q <= {(ADDR_W) {1'b0}};
      wr_ptr_q <= {(ADDR_W) {1'b0}};
    end else begin
      // Push
      if (push_i & accept_o) begin
        ram_q[wr_ptr_q] <= data_in_i;
        wr_ptr_q        <= wr_ptr_q + 1;
      end

      // Pop
      if (pop_i & valid_o) rd_ptr_q <= rd_ptr_q + 1;

      // Count up
      if ((push_i & accept_o) & ~(pop_i & valid_o)) count_q <= count_q + 1;
      // Count down
      else if (~(push_i & accept_o) & (pop_i & valid_o)) count_q <= count_q - 1;
    end

  //-------------------------------------------------------------------
  // Combinatorial
  //-------------------------------------------------------------------
  /* verilator lint_off WIDTH */
  assign valid_o    = (count_q != 0);
  assign accept_o   = (count_q != DEPTH);
  /* verilator lint_on WIDTH */

  assign data_out_o = ram_q[rd_ptr_q];

endmodule
